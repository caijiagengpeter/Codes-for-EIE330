`timescale  1ns/1ns


module  vga_pic
(
    input   wire            vga_clk     ,   
    input   wire            sys_rst_n   ,   
    input   wire    [9:0]   pix_x       ,   
    input   wire    [9:0]   pix_y       ,   

    output  reg     [15:0]  pix_data        
);

parameter   CHAR_B_H=   10'd192 ,  
            CHAR_B_V=   10'd208 ;  

parameter   CHAR_W  =   10'd256 ,   
            CHAR_H  =   10'd88  ;   

parameter   BLACK   =   16'h0000,   
            WHITE   =   16'hFFFF,   
            GOLDEN  =   16'hFEC0;   

wire    [9:0]   char_x  ;   
wire    [9:0]   char_y  ;   

reg     [255:0] char    [87:0]  ;  

assign  char_x  =   (((pix_x >= CHAR_B_H) && (pix_x < (CHAR_B_H + CHAR_W)))
                    && ((pix_y >= CHAR_B_V) && (pix_y < (CHAR_B_V + CHAR_H))))
                    ? (pix_x - CHAR_B_H) : 10'h3FF;
assign  char_y  =   (((pix_x >= CHAR_B_H) && (pix_x < (CHAR_B_H + CHAR_W)))
                    && ((pix_y >= CHAR_B_V) && (pix_y < (CHAR_B_V + CHAR_H))))
                    ? (pix_y - CHAR_B_V) : 10'h3FF;

always@(posedge vga_clk)
    begin
        char[0]  <=  256'h000000000000000000000000000000000000007FF00000000000000000000000;
        char[1]  <=  256'hFFFF00000003FFFE3FFFFF00003FFFF8000007FFFE00200000FFFFFFFFFFFF00;
        char[2]  <=  256'hFFFF80000007FFFE3FFFFF00003FFFF800001FFFFF80200000FFFFFFFFFFFF00;
        char[3]  <=  256'hFFFF80000007FFFE3FFFFF00003FFFF800007F801FF0E00000FFFFFFFFFFFF80;
        char[4]  <=  256'h0FFF80000007FFE001FFE0000000FE000000FC0003FFE00000FFC01FF801FF80;
        char[5]  <=  256'h03FF80000007FFC000FFC00000007C000003F00000FFF00001FE000FF0003F80;
        char[6]  <=  256'h01FF8000000FFF80007F8000000038000007E000007FF00001FC000FF0001F80;
        char[7]  <=  256'h01FFC000000FFF80007F800000003800000FC000003FF00001F8000FF0000F80;
        char[8]  <=  256'h01FFC000000FFF80007F800000003800000F8000001FF00001F0000FF0000FC0;
        char[9]  <=  256'h01FFC000000FFF80007F800000003800001F8000000FF00003F0000FF00007C0;
        char[10] <=  256'h01FFC000000FFF80007F800000003800003F00000007F00003E0000FF00007C0;
        char[11] <=  256'h01FFE000001FFF80007F800000003800003F00000003F00003E0000FF00003C0;
        char[12] <=  256'h01FFE000001FFF80007F800000003800007E00000003F00003C0000FF00003E0;
        char[13] <=  256'h01FFE000001FFF80007F800000003800007E00000001F00007C0000FF00001E0;
        char[14] <=  256'h01FFE000001FFF80007F80000000380000FE00000001F0000780000FF00001E0;
        char[15] <=  256'h01FFE000003FFF80007F80000000380000FC00000000F8000780000FF00000E0;
        char[16] <=  256'h01FFF000003FFF80007F80000000380000FC00000000F8000700000FF00000E0;
        char[17] <=  256'h01FFF000003FFF80007F80000000380001FC0000000078000F00000FF0000070;
        char[18] <=  256'h01FFF000003FFF80007F80000000380001FC0000000078000F00000FF0000070;
        char[19] <=  256'h01FFF000007FFF80007F80000000380001FC0000000038000600000FF0000060;
        char[20] <=  256'h01FFF800007FFF80007F80000000380001FC0000000030000000000FF0000000;
        char[21] <=  256'h01FFF800007DFF80007F80000000380001FC0000000000000000000FF0000000;
        char[22] <=  256'h01FFF800007DFF80007F80000000380001FC0000000000000000000FF0000000;
        char[23] <=  256'h01EFF80000FDFF80007F80000000380001FC0000000000000000000FF0000000;
        char[24] <=  256'h01EFF80000FDFF80007F80000000380001FE0000000000000000000FF0000000;
        char[25] <=  256'h01EFFC0000FDFF80007F80000000380001FE0000000000000000000FF0000000;
        char[26] <=  256'h01EFFC0000F9FF80007F80000000380001FE0000000000000000000FF0000000;
        char[27] <=  256'h01E7FC0000F9FF80007F80000000380000FF0000000000000000000FF0000000;
        char[28] <=  256'h01E7FC0001F9FF80007F80000000380000FF8000000000000000000FF0000000;
        char[29] <=  256'h01E7FE0001F9FF80007F80000000380000FFC000000000000000000FF0000000;
        char[30] <=  256'h01E7FE0001F1FF80007F800000003800007FE000000000000000000FF0000000;
        char[31] <=  256'h01E7FE0001F1FF80007F800000003800007FF000000000000000000FF0000000;
        char[32] <=  256'h01E3FE0003F1FF80007F800000003800003FFC00000000000000000FF0000000;
        char[33] <=  256'h01E3FE0003F1FF80007F800000003800003FFF00000000000000000FF0000000;
        char[34] <=  256'h01E3FF0003E1FF80007F800000003800001FFFC0000000000000000FF0000000;
        char[35] <=  256'h01E3FF0003E1FF80007F800000003800000FFFF0000000000000000FF0000000;
        char[36] <=  256'h01E1FF0007E1FF80007F8000000038000007FFFC000000000000000FF0000000;
        char[37] <=  256'h01E1FF0007E1FF80007F8000000038000001FFFF000000000000000FF0000000;
        char[38] <=  256'h01E1FF8007C1FF80007F8000000038000000FFFFC00000000000000FF0000000;
        char[39] <=  256'h01E1FF8007C1FF80007F80000000380000003FFFF00000000000000FF0000000;
        char[40] <=  256'h01E1FF800FC1FF80007F80000000380000001FFFFC0000000000000FF0000000;
        char[41] <=  256'h01E0FF800FC1FF80007F800000003800000007FFFF0000000000000FF0000000;
        char[42] <=  256'h01E0FF800FC1FF80007F800000003800000001FFFFC000000000000FF0000000;
        char[43] <=  256'h01E0FFC00F81FF80007F8000000038000000007FFFE000000000000FF0000000;
        char[44] <=  256'h01E0FFC00F81FF80007F8000000038000000001FFFF800000000000FF0000000;
        char[45] <=  256'h01E07FC01F81FF80007F80000000380000000007FFFC00000000000FF0000000;
        char[46] <=  256'h01E07FC01F81FF80007F80000000380000000001FFFE00000000000FF0000000;
        char[47] <=  256'h01E07FC01F01FF80007F800000003800000000007FFF00000000000FF0000000;
        char[48] <=  256'h01E07FE01F01FF80007F800000003800000000001FFF80000000000FF0000000;
        char[49] <=  256'h01E03FE03F01FF80007F8000000038000000000007FFC0000000000FF0000000;
        char[50] <=  256'h01E03FE03F01FF80007F8000000038000000000003FFE0000000000FF0000000;
        char[51] <=  256'h01E03FE03E01FF80007F8000000038000000000000FFF0000000000FF0000000;
        char[52] <=  256'h01E03FF03E01FF80007F80000000380000000000007FF8000000000FF0000000;
        char[53] <=  256'h01E03FF07E01FF80007F80000000380000000000003FF8000000000FF0000000;
        char[54] <=  256'h01E01FF07E01FF80007F80000000380000000000001FFC000000000FF0000000;
        char[55] <=  256'h01E01FF07C01FF80007F80000000380000000000000FFC000000000FF0000000;
        char[56] <=  256'h01E01FF07C01FF80007F800000003800000000000007FE000000000FF0000000;
        char[57] <=  256'h01E01FF8FC01FF80007F800000003800000000000003FE000000000FF0000000;
		  char[58] <=  256'h01E00FF8FC01FF80007F800000003800000000000003FE000000000FF0000000;
		  char[59] <=  256'h01E00FF8F801FF80007F800000003800000000000001FE000000000FF0000000;  
		  char[60] <=  256'h01E00FF8F801FF80007F800000003800000000000001FF000000000FF0000000;
        char[61] <=  256'h01E00FFCF801FF80007F800000003800000000000000FF000000000FF0000000;
	  	  char[62] <=  256'h01E00FFDF801FF80007F800000003800000000000000FF000000000FF0000000;
		  char[63] <=  256'h01E007FDF801FF80007F800000003800018000000000FF000000000FF0000000;
		  char[64] <=  256'h01E007FDF001FF80007F800000003800038000000000FF000000000FF0000000;
		  char[65] <=  256'h01E007FDF001FF80007F80000000380003C000000000FF000000000FF0000000;
		  char[66] <=  256'h01E007FFF001FF80007F80000000380003C000000000FF000000000FF0000000;
		  char[67] <=  256'h01E003FFF001FF80007F80000000380001C000000000FF000000000FF0000000;
		  char[68] <=  256'h01E003FFE001FF80007F80000000380001E000000000FF000000000FF0000000;
		  char[69] <=  256'h01E003FFE001FF80007F80000000380001E000000000FF000000000FF0000000;
		  char[70] <=  256'h01E003FFE001FF80007F80000000380001F000000000FE000000000FF0000000;
		  char[71] <=  256'h01E001FFE001FF80007F80000000380001F000000001FE000000000FF0000000;
		  char[72] <=  256'h01E001FFC001FF80003F80000000700001F000000001FE000000000FF0000000;
		  char[73] <=  256'h01E001FFC001FF80003F80000000700000F800000001FC000000000FF0000000;
        char[74] <=  256'h01E001FFC001FF80003FC0000000700000FC00000001FC000000000FF0000000;
		  char[75] <=  256'h01E001FFC001FF80003FC0000000E00000FC00000003FC000000000FF0000000;
        char[76] <=  256'h01E000FF8001FF80001FC0000000E00000FE00000003F8000000000FF0000000;
	  	  char[77] <=  256'h01E000FF8001FF80001FC0000001C00000FF00000007F0000000000FF0000000;
		  char[78] <=  256'h01E000FF8001FF80000FE0000003C00000FF00000007F0000000000FF0000000;
		  char[79] <=  256'h01E000FF8001FF80000FF00000078000007F8000000FE0000000000FF0000000;
		  char[80] <=  256'h01E0007F8001FF800007F000000F0000007FE000001FC0000000000FF0000000;
		  char[81] <=  256'h01E0007F0001FF800003F800001E0000007FF000003F80000000000FF0000000;
		  char[82] <=  256'h01E0007F0001FF800001FE00003C0000007FFC00007F00000000000FF0000000;
		  char[83] <=  256'h03F0007F0001FFC00000FF0000F80000007FFF0001FE00000000001FF8000000;
		  char[84] <=  256'h0FFC007F0007FFE000003FE007E00000007C0FE00FFC00000000003FFC000000;
		  char[85] <=  256'h7FFF803E00FFFFFE00000FFFFFC00000003801FFFFF0000000001FFFFFF80000;
		  char[86] <=  256'h7FFF803E00FFFFFE000003FFFE0000000030007FFFC0000000001FFFFFF80000;
		  char[87] <=  256'h7FFF803E00FFFFFE0000003FF00000000000000FFC00000000001FFFFFF80000;
        
    end

always@(posedge vga_clk or negedge sys_rst_n)
    if(sys_rst_n == 1'b0)
        pix_data    <= BLACK;
    else    if((((pix_x >= (CHAR_B_H - 1'b1))
                && (pix_x < (CHAR_B_H + CHAR_W -1'b1)))
                && ((pix_y >= CHAR_B_V) && (pix_y < (CHAR_B_V + CHAR_H))))
                && (char[char_y][10'd255 - char_x] == 1'b1))
        pix_data    <=  GOLDEN;
    else
        pix_data    <=  WHITE;

endmodule
